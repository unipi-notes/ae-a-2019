module sigma();