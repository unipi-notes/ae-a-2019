module alu4(output [31:0] o,
	   input [31:0] a);
   
   assign
     o = a + 4;
    
endmodule // alu
