module automata(output z, input[1:2]x, output[1:2]z);

endmodule