// Generalization of a Mealy Automata module

module name(params)
    //allocate state, newstate;

    initial
        begin
            state = //initial state
        end

    always @(posedge clock)
        begin
            state = //new state
        end

    always @(*)
endmodule