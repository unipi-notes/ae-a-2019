// State change function
module sigma(input [1:2]s, output [1:2]news, input [1:2]x);
    
endmodule